`include "interface.sv"
`include "transaction.sv"
`include "monitor.sv"
`include "driver.sv"
`include "generator.sv"
`include "environment.sv"
`include "scoreboard.sv"
`include "top.sv"